-------------------------------------------------------
-- Project : 
-- Author : juliangesche
-- Date : 2020-05-12
-- File : tb_d_flipflop.vhd
------------------------------------------------------
-- Description : 
-------------------------------------------------------
-- /
-------------------------------------------------------
