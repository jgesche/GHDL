-------------------------------------------------------
-- Project : 
-- Author : juliangesche
-- Date : 2020-05-12
-- File : d_flipflop.vhd
------------------------------------------------------
-- Description : 
-------------------------------------------------------
-- /
-------------------------------------------------------
